module Descriptor_Table (SYS_ADR, Descriptor_Line);
//Implementar memoria del sistema.
input  [63:0] SYS_ADR;
wire   [63:0] SYS_ADR;

output [95:0] Descriptor_Line;
reg   [95:0]  Descriptor_Line=0; 

endmodule 
