
module control_capa_fisica(strobe_in, ack_in, idle_in, no_response, pad_response, reception_complete, transmission_complete, ack_out, strobe_out, response, command_timeout, load_send, enable_pts_wrapper, enable_stp_wrapper, pad_state, pad_enable, reset, sd_clock);


   input           strobe_in;
   input           ack_in;
   input           idle_in;
   input           no_response;
   input [135 : 0] pad_response;
   input 	   reception_complete;
   input 	   transmission_complete;
   input 	   reset;
   input 	   sd_clock;

   output 	    ack_out;
   output 	    strobe_out;
   output [135 : 0] response;
   output 	    command_timeout;
   output 	    load_send;
   output 	    enable_pts_wrapper;
   output 	    enable_stp_wrapper;
   output 	    pad_state;
   output	    pad_enable;

   // output cmd_pin;


   wire           strobe_in;
   wire           ack_in;
   wire           idle_in;
   wire           no_response;
   wire [135 : 0] pad_response;
   wire 	   reception_complete;
   wire 	   transmission_complete;
   wire 	   reset;
   wire 	   sd_clock;

   reg  	 ack_out;
   reg 	         strobe_out;
   reg [135 : 0] response;
   reg   	 command_timeout;
   reg 	         load_send;
   reg 	         enable_pts_wrapper;
   reg 	         enable_stp_wrapper;
   reg 	         pad_state;
   reg	         pad_enable;
